** sch_path: /foss/designs/test/sweep_params/RC_sweep.sch
**.subckt RC_sweep
R1 OUT signal_in 100 m=1
C1 OUT GND .01u m=1
Vin signal_in GND pulse(0 1.8 0 1ns 1ns 5us 10us)
.save i(vin)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt





.control

*set hcopydevtype = svg
*set nolegend
*set color0=white
*set color1=black
*set color2=blue
*set color3=red



save i(out)
save v(out)

save all

let start_c = 10n
let stop_c = 100n
let delta_c = 20n

let c_act = start_c

* loop start
while c_act le stop_c

  alter c1 $&c_act
  tran 0.01n 20u
  let c_act = c_act + delta_c
end


plot tran1.v(out) tran2.v(out) tran3.v(out) tran4.v(out)
plot signal_in tran1.v(out) tran2.v(out) tran3.v(out) tran4.v(out)

.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
